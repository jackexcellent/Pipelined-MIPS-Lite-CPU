library verilog;
use verilog.vl_types.all;
entity tb_Multiplier is
end tb_Multiplier;
